zdvffdrsahera
